LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TB_MEMORI1 IS
END TB_MEMORI1;
 
ARCHITECTURE behavior OF TB_MEMORI1 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Memoria1
    PORT(
         clk : IN  std_logic;
         en : IN  std_logic;
         we : IN  std_logic;
         rst : IN  std_logic;
         addr : IN  std_logic_vector(9 downto 0);
         di : IN  std_logic_vector(15 downto 0);
         do : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal en : std_logic := '0';
   signal we : std_logic := '0';
   signal rst : std_logic := '0';
   signal addr : std_logic_vector(9 downto 0) := (others => '0');
   signal di : std_logic_vector(15 downto 0) := (others => '0');

 	--Outputs
   signal do : std_logic_vector(15 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Memoria1 PORT MAP (
          clk => clk,
          en => en,
          we => we,
          rst => rst,
          addr => addr,
          di => di,
          do => do
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
